// 240405

`default_nettype none

module SlaveSPI (
	input wire Clock,
	input wire Reset,
);
	
	

endmodule

`default_nettype wire
