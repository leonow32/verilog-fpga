`ifndef VIM828_DEFINES_VH
`define VIM828_DEFINES_VH

`define COM0 		19
`define COM1 		36
`define COM2 		18
`define COM3  		 1

`define SEG7_XFED	 2
`define SEG7_IJKN	 3

`define BIT_A		 0
`define BIT_B		 1
`define BIT_C		 2
`define BIT_D		 3
`define BIT_E		 4
`define BIT_F		 5
`define BIT_G		 6
`define BIT_H		 7
`define BIT_I		 8
`define BIT_J		 9
`define BIT_K		10
`define BIT_L		11
`define BIT_M		12
`define BIT_N		13
`define BIT_P		14

`endif