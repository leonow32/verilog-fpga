`default_nettype none
module ROM(
	input wire Clock,
	input wire Reset,
	input wire ReadEnable_i,
	input wire [11:0] Address_i,
	output reg [ 7:0] Data_o
);

	always @(posedge Clock) begin
		if(!Reset)
			Data_o <= 0;
		else if(ReadEnable_i) begin
			case(Address_i)

				// 0 4g2
				12'h000:	Data_o <= 8'h01;
				12'h001:	Data_o <= 8'hF4;
				12'h002:	Data_o <= 8'h02;
				12'h003:	Data_o <= 8'h7D;

				// 1 8.#a2
				12'h004:	Data_o <= 8'h01;
				12'h005:	Data_o <= 8'h77;
				12'h006:	Data_o <= 8'h02;
				12'h007:	Data_o <= 8'h18;

				// 2 16g2
				12'h008:	Data_o <= 8'h00;
				12'h009:	Data_o <= 8'h7D;
				12'h00A:	Data_o <= 8'h02;
				12'h00B:	Data_o <= 8'h7D;

				// 3 16-
				12'h00C:	Data_o <= 8'h00;
				12'h00D:	Data_o <= 8'h7D;
				12'h00E:	Data_o <= 8'h00;
				12'h00F:	Data_o <= 8'h00;

				// 4 16g2
				12'h010:	Data_o <= 8'h00;
				12'h011:	Data_o <= 8'h7D;
				12'h012:	Data_o <= 8'h02;
				12'h013:	Data_o <= 8'h7D;

				// 5 8c3
				12'h014:	Data_o <= 8'h00;
				12'h015:	Data_o <= 8'hFA;
				12'h016:	Data_o <= 8'h01;
				12'h017:	Data_o <= 8'hDD;

				// 6 8g2
				12'h018:	Data_o <= 8'h00;
				12'h019:	Data_o <= 8'hFA;
				12'h01A:	Data_o <= 8'h02;
				12'h01B:	Data_o <= 8'h7D;

				// 7 8f2
				12'h01C:	Data_o <= 8'h00;
				12'h01D:	Data_o <= 8'hFA;
				12'h01E:	Data_o <= 8'h02;
				12'h01F:	Data_o <= 8'hCB;

				// 8 4g2
				12'h020:	Data_o <= 8'h01;
				12'h021:	Data_o <= 8'hF4;
				12'h022:	Data_o <= 8'h02;
				12'h023:	Data_o <= 8'h7D;

				// 9 8.d3
				12'h024:	Data_o <= 8'h01;
				12'h025:	Data_o <= 8'h77;
				12'h026:	Data_o <= 8'h01;
				12'h027:	Data_o <= 8'hA9;

				// 10 16g2
				12'h028:	Data_o <= 8'h00;
				12'h029:	Data_o <= 8'h7D;
				12'h02A:	Data_o <= 8'h02;
				12'h02B:	Data_o <= 8'h7D;

				// 11 16-
				12'h02C:	Data_o <= 8'h00;
				12'h02D:	Data_o <= 8'h7D;
				12'h02E:	Data_o <= 8'h00;
				12'h02F:	Data_o <= 8'h00;

				// 12 16g2
				12'h030:	Data_o <= 8'h00;
				12'h031:	Data_o <= 8'h7D;
				12'h032:	Data_o <= 8'h02;
				12'h033:	Data_o <= 8'h7D;

				// 13 8#d3
				12'h034:	Data_o <= 8'h00;
				12'h035:	Data_o <= 8'hFA;
				12'h036:	Data_o <= 8'h01;
				12'h037:	Data_o <= 8'h91;

				// 14 8d3
				12'h038:	Data_o <= 8'h00;
				12'h039:	Data_o <= 8'hFA;
				12'h03A:	Data_o <= 8'h01;
				12'h03B:	Data_o <= 8'hA9;

				// 15 8#a2
				12'h03C:	Data_o <= 8'h00;
				12'h03D:	Data_o <= 8'hFA;
				12'h03E:	Data_o <= 8'h02;
				12'h03F:	Data_o <= 8'h18;

				// 16 8g2
				12'h040:	Data_o <= 8'h00;
				12'h041:	Data_o <= 8'hFA;
				12'h042:	Data_o <= 8'h02;
				12'h043:	Data_o <= 8'h7D;

				// 17 8d3
				12'h044:	Data_o <= 8'h00;
				12'h045:	Data_o <= 8'hFA;
				12'h046:	Data_o <= 8'h01;
				12'h047:	Data_o <= 8'hA9;

				// 18 8g3
				12'h048:	Data_o <= 8'h00;
				12'h049:	Data_o <= 8'hFA;
				12'h04A:	Data_o <= 8'h01;
				12'h04B:	Data_o <= 8'h3E;

				// 19 16g2
				12'h04C:	Data_o <= 8'h00;
				12'h04D:	Data_o <= 8'h7D;
				12'h04E:	Data_o <= 8'h02;
				12'h04F:	Data_o <= 8'h7D;

				// 20 16f2
				12'h050:	Data_o <= 8'h00;
				12'h051:	Data_o <= 8'h7D;
				12'h052:	Data_o <= 8'h02;
				12'h053:	Data_o <= 8'hCB;

				// 21 16-
				12'h054:	Data_o <= 8'h00;
				12'h055:	Data_o <= 8'h7D;
				12'h056:	Data_o <= 8'h00;
				12'h057:	Data_o <= 8'h00;

				// 22 16f2
				12'h058:	Data_o <= 8'h00;
				12'h059:	Data_o <= 8'h7D;
				12'h05A:	Data_o <= 8'h02;
				12'h05B:	Data_o <= 8'hCB;

				// 23 8d2
				12'h05C:	Data_o <= 8'h00;
				12'h05D:	Data_o <= 8'hFA;
				12'h05E:	Data_o <= 8'h03;
				12'h05F:	Data_o <= 8'h53;

				// 24 8a2
				12'h060:	Data_o <= 8'h00;
				12'h061:	Data_o <= 8'hFA;
				12'h062:	Data_o <= 8'h02;
				12'h063:	Data_o <= 8'h38;

				// 25 2g2
				12'h064:	Data_o <= 8'h03;
				12'h065:	Data_o <= 8'hE8;
				12'h066:	Data_o <= 8'h02;
				12'h067:	Data_o <= 8'h7D;

				// 26 2-
				12'h068:	Data_o <= 8'h03;
				12'h069:	Data_o <= 8'hE8;
				12'h06A:	Data_o <= 8'h00;
				12'h06B:	Data_o <= 8'h00;

				// 27 4a1
				12'h06C:	Data_o <= 8'h01;
				12'h06D:	Data_o <= 8'hF4;
				12'h06E:	Data_o <= 8'h04;
				12'h06F:	Data_o <= 8'h70;

				// 28 4a1
				12'h070:	Data_o <= 8'h01;
				12'h071:	Data_o <= 8'hF4;
				12'h072:	Data_o <= 8'h04;
				12'h073:	Data_o <= 8'h70;

				// 29 4a1
				12'h074:	Data_o <= 8'h01;
				12'h075:	Data_o <= 8'hF4;
				12'h076:	Data_o <= 8'h04;
				12'h077:	Data_o <= 8'h70;

				// 30 4f1
				12'h078:	Data_o <= 8'h01;
				12'h079:	Data_o <= 8'hF4;
				12'h07A:	Data_o <= 8'h05;
				12'h07B:	Data_o <= 8'h97;

				// 31 16c2
				12'h07C:	Data_o <= 8'h00;
				12'h07D:	Data_o <= 8'h7D;
				12'h07E:	Data_o <= 8'h03;
				12'h07F:	Data_o <= 8'hBB;

				// 32 4a1
				12'h080:	Data_o <= 8'h01;
				12'h081:	Data_o <= 8'hF4;
				12'h082:	Data_o <= 8'h04;
				12'h083:	Data_o <= 8'h70;

				// 33 4f1
				12'h084:	Data_o <= 8'h01;
				12'h085:	Data_o <= 8'hF4;
				12'h086:	Data_o <= 8'h05;
				12'h087:	Data_o <= 8'h97;

				// 34 16c2
				12'h088:	Data_o <= 8'h00;
				12'h089:	Data_o <= 8'h7D;
				12'h08A:	Data_o <= 8'h03;
				12'h08B:	Data_o <= 8'hBB;

				// 35 2a1
				12'h08C:	Data_o <= 8'h03;
				12'h08D:	Data_o <= 8'hE8;
				12'h08E:	Data_o <= 8'h04;
				12'h08F:	Data_o <= 8'h70;

				// 36 4e2
				12'h090:	Data_o <= 8'h01;
				12'h091:	Data_o <= 8'hF4;
				12'h092:	Data_o <= 8'h02;
				12'h093:	Data_o <= 8'hF6;

				// 37 4e2
				12'h094:	Data_o <= 8'h01;
				12'h095:	Data_o <= 8'hF4;
				12'h096:	Data_o <= 8'h02;
				12'h097:	Data_o <= 8'hF6;

				// 38 4e2
				12'h098:	Data_o <= 8'h01;
				12'h099:	Data_o <= 8'hF4;
				12'h09A:	Data_o <= 8'h02;
				12'h09B:	Data_o <= 8'hF6;

				// 39 4f2
				12'h09C:	Data_o <= 8'h01;
				12'h09D:	Data_o <= 8'hF4;
				12'h09E:	Data_o <= 8'h02;
				12'h09F:	Data_o <= 8'hCB;

				// 40 16c2
				12'h0A0:	Data_o <= 8'h00;
				12'h0A1:	Data_o <= 8'h7D;
				12'h0A2:	Data_o <= 8'h03;
				12'h0A3:	Data_o <= 8'hBB;

				// 41 4#g1
				12'h0A4:	Data_o <= 8'h01;
				12'h0A5:	Data_o <= 8'hF4;
				12'h0A6:	Data_o <= 8'h04;
				12'h0A7:	Data_o <= 8'hB3;

				// 42 4f1
				12'h0A8:	Data_o <= 8'h01;
				12'h0A9:	Data_o <= 8'hF4;
				12'h0AA:	Data_o <= 8'h05;
				12'h0AB:	Data_o <= 8'h97;

				// 43 16c2
				12'h0AC:	Data_o <= 8'h00;
				12'h0AD:	Data_o <= 8'h7D;
				12'h0AE:	Data_o <= 8'h03;
				12'h0AF:	Data_o <= 8'hBB;

				// 44 2a1
				12'h0B0:	Data_o <= 8'h03;
				12'h0B1:	Data_o <= 8'hE8;
				12'h0B2:	Data_o <= 8'h04;
				12'h0B3:	Data_o <= 8'h70;

				// 45 4a2
				12'h0B4:	Data_o <= 8'h01;
				12'h0B5:	Data_o <= 8'hF4;
				12'h0B6:	Data_o <= 8'h02;
				12'h0B7:	Data_o <= 8'h38;

				// 46 4a1
				12'h0B8:	Data_o <= 8'h01;
				12'h0B9:	Data_o <= 8'hF4;
				12'h0BA:	Data_o <= 8'h04;
				12'h0BB:	Data_o <= 8'h70;

				// 47 16a1
				12'h0BC:	Data_o <= 8'h00;
				12'h0BD:	Data_o <= 8'h7D;
				12'h0BE:	Data_o <= 8'h04;
				12'h0BF:	Data_o <= 8'h70;

				// 48 4a2
				12'h0C0:	Data_o <= 8'h01;
				12'h0C1:	Data_o <= 8'hF4;
				12'h0C2:	Data_o <= 8'h02;
				12'h0C3:	Data_o <= 8'h38;

				// 49 4#g2
				12'h0C4:	Data_o <= 8'h01;
				12'h0C5:	Data_o <= 8'hF4;
				12'h0C6:	Data_o <= 8'h02;
				12'h0C7:	Data_o <= 8'h59;

				// 50 16g2
				12'h0C8:	Data_o <= 8'h00;
				12'h0C9:	Data_o <= 8'h7D;
				12'h0CA:	Data_o <= 8'h02;
				12'h0CB:	Data_o <= 8'h7D;

				// 51 16#f2
				12'h0CC:	Data_o <= 8'h00;
				12'h0CD:	Data_o <= 8'h7D;
				12'h0CE:	Data_o <= 8'h02;
				12'h0CF:	Data_o <= 8'hA3;

				// 52 16f2
				12'h0D0:	Data_o <= 8'h00;
				12'h0D1:	Data_o <= 8'h7D;
				12'h0D2:	Data_o <= 8'h02;
				12'h0D3:	Data_o <= 8'hCB;

				// 53 4#f2
				12'h0D4:	Data_o <= 8'h01;
				12'h0D5:	Data_o <= 8'hF4;
				12'h0D6:	Data_o <= 8'h02;
				12'h0D7:	Data_o <= 8'hA3;

				// 54 8#a1
				12'h0D8:	Data_o <= 8'h00;
				12'h0D9:	Data_o <= 8'hFA;
				12'h0DA:	Data_o <= 8'h04;
				12'h0DB:	Data_o <= 8'h30;

				// 55 4#d2
				12'h0DC:	Data_o <= 8'h01;
				12'h0DD:	Data_o <= 8'hF4;
				12'h0DE:	Data_o <= 8'h03;
				12'h0DF:	Data_o <= 8'h23;

				// 56 4d2
				12'h0E0:	Data_o <= 8'h01;
				12'h0E1:	Data_o <= 8'hF4;
				12'h0E2:	Data_o <= 8'h03;
				12'h0E3:	Data_o <= 8'h53;

				// 57 16#c2
				12'h0E4:	Data_o <= 8'h00;
				12'h0E5:	Data_o <= 8'h7D;
				12'h0E6:	Data_o <= 8'h03;
				12'h0E7:	Data_o <= 8'h85;

				// 58 16c2
				12'h0E8:	Data_o <= 8'h00;
				12'h0E9:	Data_o <= 8'h7D;
				12'h0EA:	Data_o <= 8'h03;
				12'h0EB:	Data_o <= 8'hBB;

				// 59 16b1
				12'h0EC:	Data_o <= 8'h00;
				12'h0ED:	Data_o <= 8'h7D;
				12'h0EE:	Data_o <= 8'h03;
				12'h0EF:	Data_o <= 8'hF4;

				// 60 4c2
				12'h0F0:	Data_o <= 8'h01;
				12'h0F1:	Data_o <= 8'hF4;
				12'h0F2:	Data_o <= 8'h03;
				12'h0F3:	Data_o <= 8'hBB;

				// 61 8f1
				12'h0F4:	Data_o <= 8'h00;
				12'h0F5:	Data_o <= 8'hFA;
				12'h0F6:	Data_o <= 8'h05;
				12'h0F7:	Data_o <= 8'h97;

				// 62 4#g1
				12'h0F8:	Data_o <= 8'h01;
				12'h0F9:	Data_o <= 8'hF4;
				12'h0FA:	Data_o <= 8'h04;
				12'h0FB:	Data_o <= 8'hB3;

				// 63 4f1
				12'h0FC:	Data_o <= 8'h01;
				12'h0FD:	Data_o <= 8'hF4;
				12'h0FE:	Data_o <= 8'h05;
				12'h0FF:	Data_o <= 8'h97;

				// 64 16#g1
				12'h100:	Data_o <= 8'h00;
				12'h101:	Data_o <= 8'h7D;
				12'h102:	Data_o <= 8'h04;
				12'h103:	Data_o <= 8'hB3;

				// 65 4c2
				12'h104:	Data_o <= 8'h01;
				12'h105:	Data_o <= 8'hF4;
				12'h106:	Data_o <= 8'h03;
				12'h107:	Data_o <= 8'hBB;

				// 66 4a1
				12'h108:	Data_o <= 8'h01;
				12'h109:	Data_o <= 8'hF4;
				12'h10A:	Data_o <= 8'h04;
				12'h10B:	Data_o <= 8'h70;

				// 67 16c2
				12'h10C:	Data_o <= 8'h00;
				12'h10D:	Data_o <= 8'h7D;
				12'h10E:	Data_o <= 8'h03;
				12'h10F:	Data_o <= 8'hBB;

				// 68 2e2
				12'h110:	Data_o <= 8'h03;
				12'h111:	Data_o <= 8'hE8;
				12'h112:	Data_o <= 8'h02;
				12'h113:	Data_o <= 8'hF6;

				// 69 2-
				12'h114:	Data_o <= 8'h03;
				12'h115:	Data_o <= 8'hE8;
				12'h116:	Data_o <= 8'h00;
				12'h117:	Data_o <= 8'h00;

				// 70 8b1
				12'h118:	Data_o <= 8'h00;
				12'h119:	Data_o <= 8'hFA;
				12'h11A:	Data_o <= 8'h03;
				12'h11B:	Data_o <= 8'hF4;

				// 71 8.e2
				12'h11C:	Data_o <= 8'h01;
				12'h11D:	Data_o <= 8'h77;
				12'h11E:	Data_o <= 8'h02;
				12'h11F:	Data_o <= 8'hF6;

				// 72 16g2
				12'h120:	Data_o <= 8'h00;
				12'h121:	Data_o <= 8'h7D;
				12'h122:	Data_o <= 8'h02;
				12'h123:	Data_o <= 8'h7D;

				// 73 8#f2
				12'h124:	Data_o <= 8'h00;
				12'h125:	Data_o <= 8'hFA;
				12'h126:	Data_o <= 8'h02;
				12'h127:	Data_o <= 8'hA3;

				// 74 4e2
				12'h128:	Data_o <= 8'h01;
				12'h129:	Data_o <= 8'hF4;
				12'h12A:	Data_o <= 8'h02;
				12'h12B:	Data_o <= 8'hF6;

				// 75 8b2
				12'h12C:	Data_o <= 8'h00;
				12'h12D:	Data_o <= 8'hFA;
				12'h12E:	Data_o <= 8'h01;
				12'h12F:	Data_o <= 8'hFA;

				// 76 4.a2
				12'h130:	Data_o <= 8'h02;
				12'h131:	Data_o <= 8'hEE;
				12'h132:	Data_o <= 8'h02;
				12'h133:	Data_o <= 8'h38;

				// 77 4.#f2
				12'h134:	Data_o <= 8'h02;
				12'h135:	Data_o <= 8'hEE;
				12'h136:	Data_o <= 8'h02;
				12'h137:	Data_o <= 8'hA3;

				// 78 8.e2
				12'h138:	Data_o <= 8'h01;
				12'h139:	Data_o <= 8'h77;
				12'h13A:	Data_o <= 8'h02;
				12'h13B:	Data_o <= 8'hF6;

				// 79 16g2
				12'h13C:	Data_o <= 8'h00;
				12'h13D:	Data_o <= 8'h7D;
				12'h13E:	Data_o <= 8'h02;
				12'h13F:	Data_o <= 8'h7D;

				// 80 8#f2
				12'h140:	Data_o <= 8'h00;
				12'h141:	Data_o <= 8'hFA;
				12'h142:	Data_o <= 8'h02;
				12'h143:	Data_o <= 8'hA3;

				// 81 4d2
				12'h144:	Data_o <= 8'h01;
				12'h145:	Data_o <= 8'hF4;
				12'h146:	Data_o <= 8'h03;
				12'h147:	Data_o <= 8'h53;

				// 82 8f2
				12'h148:	Data_o <= 8'h00;
				12'h149:	Data_o <= 8'hFA;
				12'h14A:	Data_o <= 8'h02;
				12'h14B:	Data_o <= 8'hCB;

				// 83 2b1
				12'h14C:	Data_o <= 8'h03;
				12'h14D:	Data_o <= 8'hE8;
				12'h14E:	Data_o <= 8'h03;
				12'h14F:	Data_o <= 8'hF4;

				// 84 8-
				12'h150:	Data_o <= 8'h00;
				12'h151:	Data_o <= 8'hFA;
				12'h152:	Data_o <= 8'h00;
				12'h153:	Data_o <= 8'h00;

				// 85 8b1
				12'h154:	Data_o <= 8'h00;
				12'h155:	Data_o <= 8'hFA;
				12'h156:	Data_o <= 8'h03;
				12'h157:	Data_o <= 8'hF4;

				// 86 8.e2
				12'h158:	Data_o <= 8'h01;
				12'h159:	Data_o <= 8'h77;
				12'h15A:	Data_o <= 8'h02;
				12'h15B:	Data_o <= 8'hF6;

				// 87 16g2
				12'h15C:	Data_o <= 8'h00;
				12'h15D:	Data_o <= 8'h7D;
				12'h15E:	Data_o <= 8'h02;
				12'h15F:	Data_o <= 8'h7D;

				// 88 8#f2
				12'h160:	Data_o <= 8'h00;
				12'h161:	Data_o <= 8'hFA;
				12'h162:	Data_o <= 8'h02;
				12'h163:	Data_o <= 8'hA3;

				// 89 4e2
				12'h164:	Data_o <= 8'h01;
				12'h165:	Data_o <= 8'hF4;
				12'h166:	Data_o <= 8'h02;
				12'h167:	Data_o <= 8'hF6;

				// 90 8b2
				12'h168:	Data_o <= 8'h00;
				12'h169:	Data_o <= 8'hFA;
				12'h16A:	Data_o <= 8'h01;
				12'h16B:	Data_o <= 8'hFA;

				// 91 4d3
				12'h16C:	Data_o <= 8'h01;
				12'h16D:	Data_o <= 8'hF4;
				12'h16E:	Data_o <= 8'h01;
				12'h16F:	Data_o <= 8'hA9;

				// 92 8#c3
				12'h170:	Data_o <= 8'h00;
				12'h171:	Data_o <= 8'hFA;
				12'h172:	Data_o <= 8'h01;
				12'h173:	Data_o <= 8'hC2;

				// 93 4c3
				12'h174:	Data_o <= 8'h01;
				12'h175:	Data_o <= 8'hF4;
				12'h176:	Data_o <= 8'h01;
				12'h177:	Data_o <= 8'hDD;

				// 94 8#g2
				12'h178:	Data_o <= 8'h00;
				12'h179:	Data_o <= 8'hFA;
				12'h17A:	Data_o <= 8'h02;
				12'h17B:	Data_o <= 8'h59;

				// 95 8.c3
				12'h17C:	Data_o <= 8'h01;
				12'h17D:	Data_o <= 8'h77;
				12'h17E:	Data_o <= 8'h01;
				12'h17F:	Data_o <= 8'hDD;

				// 96 16b2
				12'h180:	Data_o <= 8'h00;
				12'h181:	Data_o <= 8'h7D;
				12'h182:	Data_o <= 8'h01;
				12'h183:	Data_o <= 8'hFA;

				// 97 8#a2
				12'h184:	Data_o <= 8'h00;
				12'h185:	Data_o <= 8'hFA;
				12'h186:	Data_o <= 8'h02;
				12'h187:	Data_o <= 8'h18;

				// 98 4#f2
				12'h188:	Data_o <= 8'h01;
				12'h189:	Data_o <= 8'hF4;
				12'h18A:	Data_o <= 8'h02;
				12'h18B:	Data_o <= 8'hA3;

				// 99 8g2
				12'h18C:	Data_o <= 8'h00;
				12'h18D:	Data_o <= 8'hFA;
				12'h18E:	Data_o <= 8'h02;
				12'h18F:	Data_o <= 8'h7D;

				// 100 2e2
				12'h190:	Data_o <= 8'h03;
				12'h191:	Data_o <= 8'hE8;
				12'h192:	Data_o <= 8'h02;
				12'h193:	Data_o <= 8'hF6;

				// 101 8-
				12'h194:	Data_o <= 8'h00;
				12'h195:	Data_o <= 8'hFA;
				12'h196:	Data_o <= 8'h00;
				12'h197:	Data_o <= 8'h00;

				// 102 8g2
				12'h198:	Data_o <= 8'h00;
				12'h199:	Data_o <= 8'hFA;
				12'h19A:	Data_o <= 8'h02;
				12'h19B:	Data_o <= 8'h7D;

				// 103 4b2
				12'h19C:	Data_o <= 8'h01;
				12'h19D:	Data_o <= 8'hF4;
				12'h19E:	Data_o <= 8'h01;
				12'h19F:	Data_o <= 8'hFA;

				// 104 8g2
				12'h1A0:	Data_o <= 8'h00;
				12'h1A1:	Data_o <= 8'hFA;
				12'h1A2:	Data_o <= 8'h02;
				12'h1A3:	Data_o <= 8'h7D;

				// 105 4b2
				12'h1A4:	Data_o <= 8'h01;
				12'h1A5:	Data_o <= 8'hF4;
				12'h1A6:	Data_o <= 8'h01;
				12'h1A7:	Data_o <= 8'hFA;

				// 106 8g2
				12'h1A8:	Data_o <= 8'h00;
				12'h1A9:	Data_o <= 8'hFA;
				12'h1AA:	Data_o <= 8'h02;
				12'h1AB:	Data_o <= 8'h7D;

				// 107 4c3
				12'h1AC:	Data_o <= 8'h01;
				12'h1AD:	Data_o <= 8'hF4;
				12'h1AE:	Data_o <= 8'h01;
				12'h1AF:	Data_o <= 8'hDD;

				// 108 8b2
				12'h1B0:	Data_o <= 8'h00;
				12'h1B1:	Data_o <= 8'hFA;
				12'h1B2:	Data_o <= 8'h01;
				12'h1B3:	Data_o <= 8'hFA;

				// 109 4#a2
				12'h1B4:	Data_o <= 8'h01;
				12'h1B5:	Data_o <= 8'hF4;
				12'h1B6:	Data_o <= 8'h02;
				12'h1B7:	Data_o <= 8'h18;

				// 110 8#f2
				12'h1B8:	Data_o <= 8'h00;
				12'h1B9:	Data_o <= 8'hFA;
				12'h1BA:	Data_o <= 8'h02;
				12'h1BB:	Data_o <= 8'hA3;

				// 111 8.g2
				12'h1BC:	Data_o <= 8'h01;
				12'h1BD:	Data_o <= 8'h77;
				12'h1BE:	Data_o <= 8'h02;
				12'h1BF:	Data_o <= 8'h7D;

				// 112 16b2
				12'h1C0:	Data_o <= 8'h00;
				12'h1C1:	Data_o <= 8'h7D;
				12'h1C2:	Data_o <= 8'h01;
				12'h1C3:	Data_o <= 8'hFA;

				// 113 8#a2
				12'h1C4:	Data_o <= 8'h00;
				12'h1C5:	Data_o <= 8'hFA;
				12'h1C6:	Data_o <= 8'h02;
				12'h1C7:	Data_o <= 8'h18;

				// 114 4#a1
				12'h1C8:	Data_o <= 8'h01;
				12'h1C9:	Data_o <= 8'hF4;
				12'h1CA:	Data_o <= 8'h04;
				12'h1CB:	Data_o <= 8'h30;

				// 115 2-
				12'h1CC:	Data_o <= 8'h03;
				12'h1CD:	Data_o <= 8'hE8;
				12'h1CE:	Data_o <= 8'h00;
				12'h1CF:	Data_o <= 8'h00;

				// 116 8#g1
				12'h1D0:	Data_o <= 8'h00;
				12'h1D1:	Data_o <= 8'hFA;
				12'h1D2:	Data_o <= 8'h04;
				12'h1D3:	Data_o <= 8'hB3;

				// 117 2a1
				12'h1D4:	Data_o <= 8'h03;
				12'h1D5:	Data_o <= 8'hE8;
				12'h1D6:	Data_o <= 8'h04;
				12'h1D7:	Data_o <= 8'h70;

				// 118 8b1
				12'h1D8:	Data_o <= 8'h00;
				12'h1D9:	Data_o <= 8'hFA;
				12'h1DA:	Data_o <= 8'h03;
				12'h1DB:	Data_o <= 8'hF4;

				// 119 2c2
				12'h1DC:	Data_o <= 8'h03;
				12'h1DD:	Data_o <= 8'hE8;
				12'h1DE:	Data_o <= 8'h03;
				12'h1DF:	Data_o <= 8'hBB;

				// 120 8#g1
				12'h1E0:	Data_o <= 8'h00;
				12'h1E1:	Data_o <= 8'hFA;
				12'h1E2:	Data_o <= 8'h04;
				12'h1E3:	Data_o <= 8'hB3;

				// 121 8a1
				12'h1E4:	Data_o <= 8'h00;
				12'h1E5:	Data_o <= 8'hFA;
				12'h1E6:	Data_o <= 8'h04;
				12'h1E7:	Data_o <= 8'h70;

				// 122 8b1
				12'h1E8:	Data_o <= 8'h00;
				12'h1E9:	Data_o <= 8'hFA;
				12'h1EA:	Data_o <= 8'h03;
				12'h1EB:	Data_o <= 8'hF4;

				// 123 8c2
				12'h1EC:	Data_o <= 8'h00;
				12'h1ED:	Data_o <= 8'hFA;
				12'h1EE:	Data_o <= 8'h03;
				12'h1EF:	Data_o <= 8'hBB;

				// 124 8f2
				12'h1F0:	Data_o <= 8'h00;
				12'h1F1:	Data_o <= 8'hFA;
				12'h1F2:	Data_o <= 8'h02;
				12'h1F3:	Data_o <= 8'hCB;

				// 125 8e2
				12'h1F4:	Data_o <= 8'h00;
				12'h1F5:	Data_o <= 8'hFA;
				12'h1F6:	Data_o <= 8'h02;
				12'h1F7:	Data_o <= 8'hF6;

				// 126 8a1
				12'h1F8:	Data_o <= 8'h00;
				12'h1F9:	Data_o <= 8'hFA;
				12'h1FA:	Data_o <= 8'h04;
				12'h1FB:	Data_o <= 8'h70;

				// 127 8c2
				12'h1FC:	Data_o <= 8'h00;
				12'h1FD:	Data_o <= 8'hFA;
				12'h1FE:	Data_o <= 8'h03;
				12'h1FF:	Data_o <= 8'hBB;

				// 128 8e2
				12'h200:	Data_o <= 8'h00;
				12'h201:	Data_o <= 8'hFA;
				12'h202:	Data_o <= 8'h02;
				12'h203:	Data_o <= 8'hF6;

				// 129 2#d2
				12'h204:	Data_o <= 8'h03;
				12'h205:	Data_o <= 8'hE8;
				12'h206:	Data_o <= 8'h03;
				12'h207:	Data_o <= 8'h23;

				// 130 16d2
				12'h208:	Data_o <= 8'h00;
				12'h209:	Data_o <= 8'h7D;
				12'h20A:	Data_o <= 8'h03;
				12'h20B:	Data_o <= 8'h53;

				// 131 16c2
				12'h20C:	Data_o <= 8'h00;
				12'h20D:	Data_o <= 8'h7D;
				12'h20E:	Data_o <= 8'h03;
				12'h20F:	Data_o <= 8'hBB;

				// 132 16a1
				12'h210:	Data_o <= 8'h00;
				12'h211:	Data_o <= 8'h7D;
				12'h212:	Data_o <= 8'h04;
				12'h213:	Data_o <= 8'h70;

				// 133 8g1
				12'h214:	Data_o <= 8'h00;
				12'h215:	Data_o <= 8'hFA;
				12'h216:	Data_o <= 8'h04;
				12'h217:	Data_o <= 8'hFB;

				// 134 1a1
				12'h218:	Data_o <= 8'h07;
				12'h219:	Data_o <= 8'hD0;
				12'h21A:	Data_o <= 8'h04;
				12'h21B:	Data_o <= 8'h70;

				// 135 8#g1
				12'h21C:	Data_o <= 8'h00;
				12'h21D:	Data_o <= 8'hFA;
				12'h21E:	Data_o <= 8'h04;
				12'h21F:	Data_o <= 8'hB3;

				// 136 2a1
				12'h220:	Data_o <= 8'h03;
				12'h221:	Data_o <= 8'hE8;
				12'h222:	Data_o <= 8'h04;
				12'h223:	Data_o <= 8'h70;

				// 137 8b1
				12'h224:	Data_o <= 8'h00;
				12'h225:	Data_o <= 8'hFA;
				12'h226:	Data_o <= 8'h03;
				12'h227:	Data_o <= 8'hF4;

				// 138 2c2
				12'h228:	Data_o <= 8'h03;
				12'h229:	Data_o <= 8'hE8;
				12'h22A:	Data_o <= 8'h03;
				12'h22B:	Data_o <= 8'hBB;

				// 139 8#g1
				12'h22C:	Data_o <= 8'h00;
				12'h22D:	Data_o <= 8'hFA;
				12'h22E:	Data_o <= 8'h04;
				12'h22F:	Data_o <= 8'hB3;

				// 140 8a1
				12'h230:	Data_o <= 8'h00;
				12'h231:	Data_o <= 8'hFA;
				12'h232:	Data_o <= 8'h04;
				12'h233:	Data_o <= 8'h70;

				// 141 8b1
				12'h234:	Data_o <= 8'h00;
				12'h235:	Data_o <= 8'hFA;
				12'h236:	Data_o <= 8'h03;
				12'h237:	Data_o <= 8'hF4;

				// 142 8c2
				12'h238:	Data_o <= 8'h00;
				12'h239:	Data_o <= 8'hFA;
				12'h23A:	Data_o <= 8'h03;
				12'h23B:	Data_o <= 8'hBB;

				// 143 8f2
				12'h23C:	Data_o <= 8'h00;
				12'h23D:	Data_o <= 8'hFA;
				12'h23E:	Data_o <= 8'h02;
				12'h23F:	Data_o <= 8'hCB;

				// 144 8e2
				12'h240:	Data_o <= 8'h00;
				12'h241:	Data_o <= 8'hFA;
				12'h242:	Data_o <= 8'h02;
				12'h243:	Data_o <= 8'hF6;

				// 145 8c2
				12'h244:	Data_o <= 8'h00;
				12'h245:	Data_o <= 8'hFA;
				12'h246:	Data_o <= 8'h03;
				12'h247:	Data_o <= 8'hBB;

				// 146 8e2
				12'h248:	Data_o <= 8'h00;
				12'h249:	Data_o <= 8'hFA;
				12'h24A:	Data_o <= 8'h02;
				12'h24B:	Data_o <= 8'hF6;

				// 147 8a2
				12'h24C:	Data_o <= 8'h00;
				12'h24D:	Data_o <= 8'hFA;
				12'h24E:	Data_o <= 8'h02;
				12'h24F:	Data_o <= 8'h38;

				// 148 1#g2
				12'h250:	Data_o <= 8'h07;
				12'h251:	Data_o <= 8'hD0;
				12'h252:	Data_o <= 8'h02;
				12'h253:	Data_o <= 8'h59;

				// 149 8#g1
				12'h254:	Data_o <= 8'h00;
				12'h255:	Data_o <= 8'hFA;
				12'h256:	Data_o <= 8'h04;
				12'h257:	Data_o <= 8'hB3;

				// 150 2a1
				12'h258:	Data_o <= 8'h03;
				12'h259:	Data_o <= 8'hE8;
				12'h25A:	Data_o <= 8'h04;
				12'h25B:	Data_o <= 8'h70;

				// 151 8b1
				12'h25C:	Data_o <= 8'h00;
				12'h25D:	Data_o <= 8'hFA;
				12'h25E:	Data_o <= 8'h03;
				12'h25F:	Data_o <= 8'hF4;

				// 152 2c2
				12'h260:	Data_o <= 8'h03;
				12'h261:	Data_o <= 8'hE8;
				12'h262:	Data_o <= 8'h03;
				12'h263:	Data_o <= 8'hBB;

				// 153 16#g1
				12'h264:	Data_o <= 8'h00;
				12'h265:	Data_o <= 8'h7D;
				12'h266:	Data_o <= 8'h04;
				12'h267:	Data_o <= 8'hB3;

				// 154 8a1
				12'h268:	Data_o <= 8'h00;
				12'h269:	Data_o <= 8'hFA;
				12'h26A:	Data_o <= 8'h04;
				12'h26B:	Data_o <= 8'h70;

				// 155 8b1
				12'h26C:	Data_o <= 8'h00;
				12'h26D:	Data_o <= 8'hFA;
				12'h26E:	Data_o <= 8'h03;
				12'h26F:	Data_o <= 8'hF4;

				// 156 8c2
				12'h270:	Data_o <= 8'h00;
				12'h271:	Data_o <= 8'hFA;
				12'h272:	Data_o <= 8'h03;
				12'h273:	Data_o <= 8'hBB;

				// 157 8f2
				12'h274:	Data_o <= 8'h00;
				12'h275:	Data_o <= 8'hFA;
				12'h276:	Data_o <= 8'h02;
				12'h277:	Data_o <= 8'hCB;

				// 158 8e2
				12'h278:	Data_o <= 8'h00;
				12'h279:	Data_o <= 8'hFA;
				12'h27A:	Data_o <= 8'h02;
				12'h27B:	Data_o <= 8'hF6;

				// 159 8a1
				12'h27C:	Data_o <= 8'h00;
				12'h27D:	Data_o <= 8'hFA;
				12'h27E:	Data_o <= 8'h04;
				12'h27F:	Data_o <= 8'h70;

				// 160 8c2
				12'h280:	Data_o <= 8'h00;
				12'h281:	Data_o <= 8'hFA;
				12'h282:	Data_o <= 8'h03;
				12'h283:	Data_o <= 8'hBB;

				// 161 8e2
				12'h284:	Data_o <= 8'h00;
				12'h285:	Data_o <= 8'hFA;
				12'h286:	Data_o <= 8'h02;
				12'h287:	Data_o <= 8'hF6;

				// 162 2#d2
				12'h288:	Data_o <= 8'h03;
				12'h289:	Data_o <= 8'hE8;
				12'h28A:	Data_o <= 8'h03;
				12'h28B:	Data_o <= 8'h23;

				// 163 8d2
				12'h28C:	Data_o <= 8'h00;
				12'h28D:	Data_o <= 8'hFA;
				12'h28E:	Data_o <= 8'h03;
				12'h28F:	Data_o <= 8'h53;

				// 164 16c2
				12'h290:	Data_o <= 8'h00;
				12'h291:	Data_o <= 8'h7D;
				12'h292:	Data_o <= 8'h03;
				12'h293:	Data_o <= 8'hBB;

				// 165 16a1
				12'h294:	Data_o <= 8'h00;
				12'h295:	Data_o <= 8'h7D;
				12'h296:	Data_o <= 8'h04;
				12'h297:	Data_o <= 8'h70;

				// 166 2-
				12'h298:	Data_o <= 8'h03;
				12'h299:	Data_o <= 8'hE8;
				12'h29A:	Data_o <= 8'h00;
				12'h29B:	Data_o <= 8'h00;

				// 167 8#c1
				12'h29C:	Data_o <= 8'h00;
				12'h29D:	Data_o <= 8'hFA;
				12'h29E:	Data_o <= 8'h07;
				12'h29F:	Data_o <= 8'h0B;

				// 168 8#c1
				12'h2A0:	Data_o <= 8'h00;
				12'h2A1:	Data_o <= 8'hFA;
				12'h2A2:	Data_o <= 8'h07;
				12'h2A3:	Data_o <= 8'h0B;

				// 169 16#c1
				12'h2A4:	Data_o <= 8'h00;
				12'h2A5:	Data_o <= 8'h7D;
				12'h2A6:	Data_o <= 8'h07;
				12'h2A7:	Data_o <= 8'h0B;

				// 170 2#f1
				12'h2A8:	Data_o <= 8'h03;
				12'h2A9:	Data_o <= 8'hE8;
				12'h2AA:	Data_o <= 8'h05;
				12'h2AB:	Data_o <= 8'h47;

				// 171 2#c2
				12'h2AC:	Data_o <= 8'h03;
				12'h2AD:	Data_o <= 8'hE8;
				12'h2AE:	Data_o <= 8'h03;
				12'h2AF:	Data_o <= 8'h85;

				// 172 8b1
				12'h2B0:	Data_o <= 8'h00;
				12'h2B1:	Data_o <= 8'hFA;
				12'h2B2:	Data_o <= 8'h03;
				12'h2B3:	Data_o <= 8'hF4;

				// 173 16#a1
				12'h2B4:	Data_o <= 8'h00;
				12'h2B5:	Data_o <= 8'h7D;
				12'h2B6:	Data_o <= 8'h04;
				12'h2B7:	Data_o <= 8'h30;

				// 174 8#g1
				12'h2B8:	Data_o <= 8'h00;
				12'h2B9:	Data_o <= 8'hFA;
				12'h2BA:	Data_o <= 8'h04;
				12'h2BB:	Data_o <= 8'hB3;

				// 175 2#f2
				12'h2BC:	Data_o <= 8'h03;
				12'h2BD:	Data_o <= 8'hE8;
				12'h2BE:	Data_o <= 8'h02;
				12'h2BF:	Data_o <= 8'hA3;

				// 176 4#c2
				12'h2C0:	Data_o <= 8'h01;
				12'h2C1:	Data_o <= 8'hF4;
				12'h2C2:	Data_o <= 8'h03;
				12'h2C3:	Data_o <= 8'h85;

				// 177 8b1
				12'h2C4:	Data_o <= 8'h00;
				12'h2C5:	Data_o <= 8'hFA;
				12'h2C6:	Data_o <= 8'h03;
				12'h2C7:	Data_o <= 8'hF4;

				// 178 16#a1
				12'h2C8:	Data_o <= 8'h00;
				12'h2C9:	Data_o <= 8'h7D;
				12'h2CA:	Data_o <= 8'h04;
				12'h2CB:	Data_o <= 8'h30;

				// 179 8#g1
				12'h2CC:	Data_o <= 8'h00;
				12'h2CD:	Data_o <= 8'hFA;
				12'h2CE:	Data_o <= 8'h04;
				12'h2CF:	Data_o <= 8'hB3;

				// 180 2#f2
				12'h2D0:	Data_o <= 8'h03;
				12'h2D1:	Data_o <= 8'hE8;
				12'h2D2:	Data_o <= 8'h02;
				12'h2D3:	Data_o <= 8'hA3;

				// 181 4#c2
				12'h2D4:	Data_o <= 8'h01;
				12'h2D5:	Data_o <= 8'hF4;
				12'h2D6:	Data_o <= 8'h03;
				12'h2D7:	Data_o <= 8'h85;

				// 182 8b1
				12'h2D8:	Data_o <= 8'h00;
				12'h2D9:	Data_o <= 8'hFA;
				12'h2DA:	Data_o <= 8'h03;
				12'h2DB:	Data_o <= 8'hF4;

				// 183 16#a1
				12'h2DC:	Data_o <= 8'h00;
				12'h2DD:	Data_o <= 8'h7D;
				12'h2DE:	Data_o <= 8'h04;
				12'h2DF:	Data_o <= 8'h30;

				// 184 8b1
				12'h2E0:	Data_o <= 8'h00;
				12'h2E1:	Data_o <= 8'hFA;
				12'h2E2:	Data_o <= 8'h03;
				12'h2E3:	Data_o <= 8'hF4;

				// 185 2#g1
				12'h2E4:	Data_o <= 8'h03;
				12'h2E5:	Data_o <= 8'hE8;
				12'h2E6:	Data_o <= 8'h04;
				12'h2E7:	Data_o <= 8'hB3;

				// 186 8#c1
				12'h2E8:	Data_o <= 8'h00;
				12'h2E9:	Data_o <= 8'hFA;
				12'h2EA:	Data_o <= 8'h07;
				12'h2EB:	Data_o <= 8'h0B;

				// 187 8#c1
				12'h2EC:	Data_o <= 8'h00;
				12'h2ED:	Data_o <= 8'hFA;
				12'h2EE:	Data_o <= 8'h07;
				12'h2EF:	Data_o <= 8'h0B;

				// 188 16#c1
				12'h2F0:	Data_o <= 8'h00;
				12'h2F1:	Data_o <= 8'h7D;
				12'h2F2:	Data_o <= 8'h07;
				12'h2F3:	Data_o <= 8'h0B;

				// 189 2#f1
				12'h2F4:	Data_o <= 8'h03;
				12'h2F5:	Data_o <= 8'hE8;
				12'h2F6:	Data_o <= 8'h05;
				12'h2F7:	Data_o <= 8'h47;

				// 190 2#c2
				12'h2F8:	Data_o <= 8'h03;
				12'h2F9:	Data_o <= 8'hE8;
				12'h2FA:	Data_o <= 8'h03;
				12'h2FB:	Data_o <= 8'h85;

				// 191 8b1
				12'h2FC:	Data_o <= 8'h00;
				12'h2FD:	Data_o <= 8'hFA;
				12'h2FE:	Data_o <= 8'h03;
				12'h2FF:	Data_o <= 8'hF4;

				// 192 16#a1
				12'h300:	Data_o <= 8'h00;
				12'h301:	Data_o <= 8'h7D;
				12'h302:	Data_o <= 8'h04;
				12'h303:	Data_o <= 8'h30;

				// 193 8#g1
				12'h304:	Data_o <= 8'h00;
				12'h305:	Data_o <= 8'hFA;
				12'h306:	Data_o <= 8'h04;
				12'h307:	Data_o <= 8'hB3;

				// 194 2#f2
				12'h308:	Data_o <= 8'h03;
				12'h309:	Data_o <= 8'hE8;
				12'h30A:	Data_o <= 8'h02;
				12'h30B:	Data_o <= 8'hA3;

				// 195 4#c2
				12'h30C:	Data_o <= 8'h01;
				12'h30D:	Data_o <= 8'hF4;
				12'h30E:	Data_o <= 8'h03;
				12'h30F:	Data_o <= 8'h85;

				// 196 8b1
				12'h310:	Data_o <= 8'h00;
				12'h311:	Data_o <= 8'hFA;
				12'h312:	Data_o <= 8'h03;
				12'h313:	Data_o <= 8'hF4;

				// 197 16#a1
				12'h314:	Data_o <= 8'h00;
				12'h315:	Data_o <= 8'h7D;
				12'h316:	Data_o <= 8'h04;
				12'h317:	Data_o <= 8'h30;

				// 198 8#g1
				12'h318:	Data_o <= 8'h00;
				12'h319:	Data_o <= 8'hFA;
				12'h31A:	Data_o <= 8'h04;
				12'h31B:	Data_o <= 8'hB3;

				// 199 2#f2
				12'h31C:	Data_o <= 8'h03;
				12'h31D:	Data_o <= 8'hE8;
				12'h31E:	Data_o <= 8'h02;
				12'h31F:	Data_o <= 8'hA3;

				// 200 4#c2
				12'h320:	Data_o <= 8'h01;
				12'h321:	Data_o <= 8'hF4;
				12'h322:	Data_o <= 8'h03;
				12'h323:	Data_o <= 8'h85;

				// 201 8b1
				12'h324:	Data_o <= 8'h00;
				12'h325:	Data_o <= 8'hFA;
				12'h326:	Data_o <= 8'h03;
				12'h327:	Data_o <= 8'hF4;

				// 202 16#a1
				12'h328:	Data_o <= 8'h00;
				12'h329:	Data_o <= 8'h7D;
				12'h32A:	Data_o <= 8'h04;
				12'h32B:	Data_o <= 8'h30;

				// 203 8b1
				12'h32C:	Data_o <= 8'h00;
				12'h32D:	Data_o <= 8'hFA;
				12'h32E:	Data_o <= 8'h03;
				12'h32F:	Data_o <= 8'hF4;

				// 204 2#g1
				12'h330:	Data_o <= 8'h03;
				12'h331:	Data_o <= 8'hE8;
				12'h332:	Data_o <= 8'h04;
				12'h333:	Data_o <= 8'hB3;

				// 205 4#c1
				12'h334:	Data_o <= 8'h01;
				12'h335:	Data_o <= 8'hF4;
				12'h336:	Data_o <= 8'h07;
				12'h337:	Data_o <= 8'h0B;

				// 206 16#c1
				12'h338:	Data_o <= 8'h00;
				12'h339:	Data_o <= 8'h7D;
				12'h33A:	Data_o <= 8'h07;
				12'h33B:	Data_o <= 8'h0B;

				// 207 2#d1
				12'h33C:	Data_o <= 8'h03;
				12'h33D:	Data_o <= 8'hE8;
				12'h33E:	Data_o <= 8'h06;
				12'h33F:	Data_o <= 8'h47;

				// 208 8#c2
				12'h340:	Data_o <= 8'h00;
				12'h341:	Data_o <= 8'hFA;
				12'h342:	Data_o <= 8'h03;
				12'h343:	Data_o <= 8'h85;

				// 209 8b1
				12'h344:	Data_o <= 8'h00;
				12'h345:	Data_o <= 8'hFA;
				12'h346:	Data_o <= 8'h03;
				12'h347:	Data_o <= 8'hF4;

				// 210 8#a1
				12'h348:	Data_o <= 8'h00;
				12'h349:	Data_o <= 8'hFA;
				12'h34A:	Data_o <= 8'h04;
				12'h34B:	Data_o <= 8'h30;

				// 211 8#g1
				12'h34C:	Data_o <= 8'h00;
				12'h34D:	Data_o <= 8'hFA;
				12'h34E:	Data_o <= 8'h04;
				12'h34F:	Data_o <= 8'hB3;

				// 212 8#f1
				12'h350:	Data_o <= 8'h00;
				12'h351:	Data_o <= 8'hFA;
				12'h352:	Data_o <= 8'h05;
				12'h353:	Data_o <= 8'h47;

				// 213 16#f1
				12'h354:	Data_o <= 8'h00;
				12'h355:	Data_o <= 8'h7D;
				12'h356:	Data_o <= 8'h05;
				12'h357:	Data_o <= 8'h47;

				// 214 8#g1
				12'h358:	Data_o <= 8'h00;
				12'h359:	Data_o <= 8'hFA;
				12'h35A:	Data_o <= 8'h04;
				12'h35B:	Data_o <= 8'hB3;

				// 215 16#a1
				12'h35C:	Data_o <= 8'h00;
				12'h35D:	Data_o <= 8'h7D;
				12'h35E:	Data_o <= 8'h04;
				12'h35F:	Data_o <= 8'h30;

				// 216 4#g1
				12'h360:	Data_o <= 8'h01;
				12'h361:	Data_o <= 8'hF4;
				12'h362:	Data_o <= 8'h04;
				12'h363:	Data_o <= 8'hB3;

				// 217 2-
				12'h364:	Data_o <= 8'h03;
				12'h365:	Data_o <= 8'hE8;
				12'h366:	Data_o <= 8'h00;
				12'h367:	Data_o <= 8'h00;

				// 218 4-
				12'h368:	Data_o <= 8'h01;
				12'h369:	Data_o <= 8'hF4;
				12'h36A:	Data_o <= 8'h00;
				12'h36B:	Data_o <= 8'h00;

				// 219 8-
				12'h36C:	Data_o <= 8'h00;
				12'h36D:	Data_o <= 8'hFA;
				12'h36E:	Data_o <= 8'h00;
				12'h36F:	Data_o <= 8'h00;

				// 220 16b2
				12'h370:	Data_o <= 8'h00;
				12'h371:	Data_o <= 8'h7D;
				12'h372:	Data_o <= 8'h01;
				12'h373:	Data_o <= 8'hFA;

				// 221 16a2
				12'h374:	Data_o <= 8'h00;
				12'h375:	Data_o <= 8'h7D;
				12'h376:	Data_o <= 8'h02;
				12'h377:	Data_o <= 8'h38;

				// 222 4b2
				12'h378:	Data_o <= 8'h01;
				12'h379:	Data_o <= 8'hF4;
				12'h37A:	Data_o <= 8'h01;
				12'h37B:	Data_o <= 8'hFA;

				// 223 4e2
				12'h37C:	Data_o <= 8'h01;
				12'h37D:	Data_o <= 8'hF4;
				12'h37E:	Data_o <= 8'h02;
				12'h37F:	Data_o <= 8'hF6;

				// 224 4-
				12'h380:	Data_o <= 8'h01;
				12'h381:	Data_o <= 8'hF4;
				12'h382:	Data_o <= 8'h00;
				12'h383:	Data_o <= 8'h00;

				// 225 8-
				12'h384:	Data_o <= 8'h00;
				12'h385:	Data_o <= 8'hFA;
				12'h386:	Data_o <= 8'h00;
				12'h387:	Data_o <= 8'h00;

				// 226 16c3
				12'h388:	Data_o <= 8'h00;
				12'h389:	Data_o <= 8'h7D;
				12'h38A:	Data_o <= 8'h01;
				12'h38B:	Data_o <= 8'hDD;

				// 227 16b2
				12'h38C:	Data_o <= 8'h00;
				12'h38D:	Data_o <= 8'h7D;
				12'h38E:	Data_o <= 8'h01;
				12'h38F:	Data_o <= 8'hFA;

				// 228 8c3
				12'h390:	Data_o <= 8'h00;
				12'h391:	Data_o <= 8'hFA;
				12'h392:	Data_o <= 8'h01;
				12'h393:	Data_o <= 8'hDD;

				// 229 8b2
				12'h394:	Data_o <= 8'h00;
				12'h395:	Data_o <= 8'hFA;
				12'h396:	Data_o <= 8'h01;
				12'h397:	Data_o <= 8'hFA;

				// 230 4a2
				12'h398:	Data_o <= 8'h01;
				12'h399:	Data_o <= 8'hF4;
				12'h39A:	Data_o <= 8'h02;
				12'h39B:	Data_o <= 8'h38;

				// 231 4-
				12'h39C:	Data_o <= 8'h01;
				12'h39D:	Data_o <= 8'hF4;
				12'h39E:	Data_o <= 8'h00;
				12'h39F:	Data_o <= 8'h00;

				// 232 8-
				12'h3A0:	Data_o <= 8'h00;
				12'h3A1:	Data_o <= 8'hFA;
				12'h3A2:	Data_o <= 8'h00;
				12'h3A3:	Data_o <= 8'h00;

				// 233 16c3
				12'h3A4:	Data_o <= 8'h00;
				12'h3A5:	Data_o <= 8'h7D;
				12'h3A6:	Data_o <= 8'h01;
				12'h3A7:	Data_o <= 8'hDD;

				// 234 16b2
				12'h3A8:	Data_o <= 8'h00;
				12'h3A9:	Data_o <= 8'h7D;
				12'h3AA:	Data_o <= 8'h01;
				12'h3AB:	Data_o <= 8'hFA;

				// 235 4c3
				12'h3AC:	Data_o <= 8'h01;
				12'h3AD:	Data_o <= 8'hF4;
				12'h3AE:	Data_o <= 8'h01;
				12'h3AF:	Data_o <= 8'hDD;

				// 236 4e2
				12'h3B0:	Data_o <= 8'h01;
				12'h3B1:	Data_o <= 8'hF4;
				12'h3B2:	Data_o <= 8'h02;
				12'h3B3:	Data_o <= 8'hF6;

				// 237 4-
				12'h3B4:	Data_o <= 8'h01;
				12'h3B5:	Data_o <= 8'hF4;
				12'h3B6:	Data_o <= 8'h00;
				12'h3B7:	Data_o <= 8'h00;

				// 238 8-
				12'h3B8:	Data_o <= 8'h00;
				12'h3B9:	Data_o <= 8'hFA;
				12'h3BA:	Data_o <= 8'h00;
				12'h3BB:	Data_o <= 8'h00;

				// 239 16a2
				12'h3BC:	Data_o <= 8'h00;
				12'h3BD:	Data_o <= 8'h7D;
				12'h3BE:	Data_o <= 8'h02;
				12'h3BF:	Data_o <= 8'h38;

				// 240 16g2
				12'h3C0:	Data_o <= 8'h00;
				12'h3C1:	Data_o <= 8'h7D;
				12'h3C2:	Data_o <= 8'h02;
				12'h3C3:	Data_o <= 8'h7D;

				// 241 8a2
				12'h3C4:	Data_o <= 8'h00;
				12'h3C5:	Data_o <= 8'hFA;
				12'h3C6:	Data_o <= 8'h02;
				12'h3C7:	Data_o <= 8'h38;

				// 242 8g2
				12'h3C8:	Data_o <= 8'h00;
				12'h3C9:	Data_o <= 8'hFA;
				12'h3CA:	Data_o <= 8'h02;
				12'h3CB:	Data_o <= 8'h7D;

				// 243 8#f2
				12'h3CC:	Data_o <= 8'h00;
				12'h3CD:	Data_o <= 8'hFA;
				12'h3CE:	Data_o <= 8'h02;
				12'h3CF:	Data_o <= 8'hA3;

				// 244 8a2
				12'h3D0:	Data_o <= 8'h00;
				12'h3D1:	Data_o <= 8'hFA;
				12'h3D2:	Data_o <= 8'h02;
				12'h3D3:	Data_o <= 8'h38;

				// 245 4g2
				12'h3D4:	Data_o <= 8'h01;
				12'h3D5:	Data_o <= 8'hF4;
				12'h3D6:	Data_o <= 8'h02;
				12'h3D7:	Data_o <= 8'h7D;

				// 246 8-
				12'h3D8:	Data_o <= 8'h00;
				12'h3D9:	Data_o <= 8'hFA;
				12'h3DA:	Data_o <= 8'h00;
				12'h3DB:	Data_o <= 8'h00;

				// 247 16#f2
				12'h3DC:	Data_o <= 8'h00;
				12'h3DD:	Data_o <= 8'h7D;
				12'h3DE:	Data_o <= 8'h02;
				12'h3DF:	Data_o <= 8'hA3;

				// 248 16g2
				12'h3E0:	Data_o <= 8'h00;
				12'h3E1:	Data_o <= 8'h7D;
				12'h3E2:	Data_o <= 8'h02;
				12'h3E3:	Data_o <= 8'h7D;

				// 249 4a2
				12'h3E4:	Data_o <= 8'h01;
				12'h3E5:	Data_o <= 8'hF4;
				12'h3E6:	Data_o <= 8'h02;
				12'h3E7:	Data_o <= 8'h38;

				// 250 8-
				12'h3E8:	Data_o <= 8'h00;
				12'h3E9:	Data_o <= 8'hFA;
				12'h3EA:	Data_o <= 8'h00;
				12'h3EB:	Data_o <= 8'h00;

				// 251 16g2
				12'h3EC:	Data_o <= 8'h00;
				12'h3ED:	Data_o <= 8'h7D;
				12'h3EE:	Data_o <= 8'h02;
				12'h3EF:	Data_o <= 8'h7D;

				// 252 16a2
				12'h3F0:	Data_o <= 8'h00;
				12'h3F1:	Data_o <= 8'h7D;
				12'h3F2:	Data_o <= 8'h02;
				12'h3F3:	Data_o <= 8'h38;

				// 253 8b2
				12'h3F4:	Data_o <= 8'h00;
				12'h3F5:	Data_o <= 8'hFA;
				12'h3F6:	Data_o <= 8'h01;
				12'h3F7:	Data_o <= 8'hFA;

				// 254 8a2
				12'h3F8:	Data_o <= 8'h00;
				12'h3F9:	Data_o <= 8'hFA;
				12'h3FA:	Data_o <= 8'h02;
				12'h3FB:	Data_o <= 8'h38;

				// 255 8g2
				12'h3FC:	Data_o <= 8'h00;
				12'h3FD:	Data_o <= 8'hFA;
				12'h3FE:	Data_o <= 8'h02;
				12'h3FF:	Data_o <= 8'h7D;

				// 256 8#f2
				12'h400:	Data_o <= 8'h00;
				12'h401:	Data_o <= 8'hFA;
				12'h402:	Data_o <= 8'h02;
				12'h403:	Data_o <= 8'hA3;

				// 257 4e2
				12'h404:	Data_o <= 8'h01;
				12'h405:	Data_o <= 8'hF4;
				12'h406:	Data_o <= 8'h02;
				12'h407:	Data_o <= 8'hF6;

				// 258 4c3
				12'h408:	Data_o <= 8'h01;
				12'h409:	Data_o <= 8'hF4;
				12'h40A:	Data_o <= 8'h01;
				12'h40B:	Data_o <= 8'hDD;

				// 259 2b2
				12'h40C:	Data_o <= 8'h03;
				12'h40D:	Data_o <= 8'hE8;
				12'h40E:	Data_o <= 8'h01;
				12'h40F:	Data_o <= 8'hFA;

				// 260 4-
				12'h410:	Data_o <= 8'h01;
				12'h411:	Data_o <= 8'hF4;
				12'h412:	Data_o <= 8'h00;
				12'h413:	Data_o <= 8'h00;

				// 261 16b2
				12'h414:	Data_o <= 8'h00;
				12'h415:	Data_o <= 8'h7D;
				12'h416:	Data_o <= 8'h01;
				12'h417:	Data_o <= 8'hFA;

				// 262 16c3
				12'h418:	Data_o <= 8'h00;
				12'h419:	Data_o <= 8'h7D;
				12'h41A:	Data_o <= 8'h01;
				12'h41B:	Data_o <= 8'hDD;

				// 263 16b2
				12'h41C:	Data_o <= 8'h00;
				12'h41D:	Data_o <= 8'h7D;
				12'h41E:	Data_o <= 8'h01;
				12'h41F:	Data_o <= 8'hFA;

				// 264 16a2
				12'h420:	Data_o <= 8'h00;
				12'h421:	Data_o <= 8'h7D;
				12'h422:	Data_o <= 8'h02;
				12'h423:	Data_o <= 8'h38;

				// 265 1b2
				12'h424:	Data_o <= 8'h07;
				12'h425:	Data_o <= 8'hD0;
				12'h426:	Data_o <= 8'h01;
				12'h427:	Data_o <= 8'hFA;

				// 266 2-
				12'h428:	Data_o <= 8'h03;
				12'h429:	Data_o <= 8'hE8;
				12'h42A:	Data_o <= 8'h00;
				12'h42B:	Data_o <= 8'h00;

				// 267 4e1
				12'h42C:	Data_o <= 8'h01;
				12'h42D:	Data_o <= 8'hF4;
				12'h42E:	Data_o <= 8'h05;
				12'h42F:	Data_o <= 8'hEC;

				// 268 4a1
				12'h430:	Data_o <= 8'h01;
				12'h431:	Data_o <= 8'hF4;
				12'h432:	Data_o <= 8'h04;
				12'h433:	Data_o <= 8'h70;

				// 269 4e1
				12'h434:	Data_o <= 8'h01;
				12'h435:	Data_o <= 8'hF4;
				12'h436:	Data_o <= 8'h05;
				12'h437:	Data_o <= 8'hEC;

				// 270 4g1
				12'h438:	Data_o <= 8'h01;
				12'h439:	Data_o <= 8'hF4;
				12'h43A:	Data_o <= 8'h04;
				12'h43B:	Data_o <= 8'hFB;

				// 271 8f1
				12'h43C:	Data_o <= 8'h00;
				12'h43D:	Data_o <= 8'hFA;
				12'h43E:	Data_o <= 8'h05;
				12'h43F:	Data_o <= 8'h97;

				// 272 2f1
				12'h440:	Data_o <= 8'h03;
				12'h441:	Data_o <= 8'hE8;
				12'h442:	Data_o <= 8'h05;
				12'h443:	Data_o <= 8'h97;

				// 273 4d1
				12'h444:	Data_o <= 8'h01;
				12'h445:	Data_o <= 8'hF4;
				12'h446:	Data_o <= 8'h06;
				12'h447:	Data_o <= 8'hA6;

				// 274 4g1
				12'h448:	Data_o <= 8'h01;
				12'h449:	Data_o <= 8'hF4;
				12'h44A:	Data_o <= 8'h04;
				12'h44B:	Data_o <= 8'hFB;

				// 275 8d1
				12'h44C:	Data_o <= 8'h00;
				12'h44D:	Data_o <= 8'hFA;
				12'h44E:	Data_o <= 8'h06;
				12'h44F:	Data_o <= 8'hA6;

				// 276 1e1
				12'h450:	Data_o <= 8'h07;
				12'h451:	Data_o <= 8'hD0;
				12'h452:	Data_o <= 8'h05;
				12'h453:	Data_o <= 8'hEC;

				// 277 4e1
				12'h454:	Data_o <= 8'h01;
				12'h455:	Data_o <= 8'hF4;
				12'h456:	Data_o <= 8'h05;
				12'h457:	Data_o <= 8'hEC;

				// 278 4a1
				12'h458:	Data_o <= 8'h01;
				12'h459:	Data_o <= 8'hF4;
				12'h45A:	Data_o <= 8'h04;
				12'h45B:	Data_o <= 8'h70;

				// 279 4e1
				12'h45C:	Data_o <= 8'h01;
				12'h45D:	Data_o <= 8'hF4;
				12'h45E:	Data_o <= 8'h05;
				12'h45F:	Data_o <= 8'hEC;

				// 280 4g1
				12'h460:	Data_o <= 8'h01;
				12'h461:	Data_o <= 8'hF4;
				12'h462:	Data_o <= 8'h04;
				12'h463:	Data_o <= 8'hFB;

				// 281 8f1
				12'h464:	Data_o <= 8'h00;
				12'h465:	Data_o <= 8'hFA;
				12'h466:	Data_o <= 8'h05;
				12'h467:	Data_o <= 8'h97;

				// 282 2f1
				12'h468:	Data_o <= 8'h03;
				12'h469:	Data_o <= 8'hE8;
				12'h46A:	Data_o <= 8'h05;
				12'h46B:	Data_o <= 8'h97;

				// 283 4d1
				12'h46C:	Data_o <= 8'h01;
				12'h46D:	Data_o <= 8'hF4;
				12'h46E:	Data_o <= 8'h06;
				12'h46F:	Data_o <= 8'hA6;

				// 284 4g1
				12'h470:	Data_o <= 8'h01;
				12'h471:	Data_o <= 8'hF4;
				12'h472:	Data_o <= 8'h04;
				12'h473:	Data_o <= 8'hFB;

				// 285 8d1
				12'h474:	Data_o <= 8'h00;
				12'h475:	Data_o <= 8'hFA;
				12'h476:	Data_o <= 8'h06;
				12'h477:	Data_o <= 8'hA6;

				// 286 1e1
				12'h478:	Data_o <= 8'h07;
				12'h479:	Data_o <= 8'hD0;
				12'h47A:	Data_o <= 8'h05;
				12'h47B:	Data_o <= 8'hEC;

				// 287 4e1
				12'h47C:	Data_o <= 8'h01;
				12'h47D:	Data_o <= 8'hF4;
				12'h47E:	Data_o <= 8'h05;
				12'h47F:	Data_o <= 8'hEC;

				// 288 4a1
				12'h480:	Data_o <= 8'h01;
				12'h481:	Data_o <= 8'hF4;
				12'h482:	Data_o <= 8'h04;
				12'h483:	Data_o <= 8'h70;

				// 289 4c2
				12'h484:	Data_o <= 8'h01;
				12'h485:	Data_o <= 8'hF4;
				12'h486:	Data_o <= 8'h03;
				12'h487:	Data_o <= 8'hBB;

				// 290 4e2
				12'h488:	Data_o <= 8'h01;
				12'h489:	Data_o <= 8'hF4;
				12'h48A:	Data_o <= 8'h02;
				12'h48B:	Data_o <= 8'hF6;

				// 291 8d2
				12'h48C:	Data_o <= 8'h00;
				12'h48D:	Data_o <= 8'hFA;
				12'h48E:	Data_o <= 8'h03;
				12'h48F:	Data_o <= 8'h53;

				// 292 2d2
				12'h490:	Data_o <= 8'h03;
				12'h491:	Data_o <= 8'hE8;
				12'h492:	Data_o <= 8'h03;
				12'h493:	Data_o <= 8'h53;

				// 293 4d2
				12'h494:	Data_o <= 8'h01;
				12'h495:	Data_o <= 8'hF4;
				12'h496:	Data_o <= 8'h03;
				12'h497:	Data_o <= 8'h53;

				// 294 4g2
				12'h498:	Data_o <= 8'h01;
				12'h499:	Data_o <= 8'hF4;
				12'h49A:	Data_o <= 8'h02;
				12'h49B:	Data_o <= 8'h7D;

				// 295 8d2
				12'h49C:	Data_o <= 8'h00;
				12'h49D:	Data_o <= 8'hFA;
				12'h49E:	Data_o <= 8'h03;
				12'h49F:	Data_o <= 8'h53;

				// 296 1e2
				12'h4A0:	Data_o <= 8'h07;
				12'h4A1:	Data_o <= 8'hD0;
				12'h4A2:	Data_o <= 8'h02;
				12'h4A3:	Data_o <= 8'hF6;

				// 297 4e2
				12'h4A4:	Data_o <= 8'h01;
				12'h4A5:	Data_o <= 8'hF4;
				12'h4A6:	Data_o <= 8'h02;
				12'h4A7:	Data_o <= 8'hF6;

				// 298 1a2
				12'h4A8:	Data_o <= 8'h07;
				12'h4A9:	Data_o <= 8'hD0;
				12'h4AA:	Data_o <= 8'h02;
				12'h4AB:	Data_o <= 8'h38;

				// 299 8g2
				12'h4AC:	Data_o <= 8'h00;
				12'h4AD:	Data_o <= 8'hFA;
				12'h4AE:	Data_o <= 8'h02;
				12'h4AF:	Data_o <= 8'h7D;

				// 300 8f2
				12'h4B0:	Data_o <= 8'h00;
				12'h4B1:	Data_o <= 8'hFA;
				12'h4B2:	Data_o <= 8'h02;
				12'h4B3:	Data_o <= 8'hCB;

				// 301 8e2
				12'h4B4:	Data_o <= 8'h00;
				12'h4B5:	Data_o <= 8'hFA;
				12'h4B6:	Data_o <= 8'h02;
				12'h4B7:	Data_o <= 8'hF6;

				// 302 8d2
				12'h4B8:	Data_o <= 8'h00;
				12'h4B9:	Data_o <= 8'hFA;
				12'h4BA:	Data_o <= 8'h03;
				12'h4BB:	Data_o <= 8'h53;

				// 303 8c2
				12'h4BC:	Data_o <= 8'h00;
				12'h4BD:	Data_o <= 8'hFA;
				12'h4BE:	Data_o <= 8'h03;
				12'h4BF:	Data_o <= 8'hBB;

				// 304 8b1
				12'h4C0:	Data_o <= 8'h00;
				12'h4C1:	Data_o <= 8'hFA;
				12'h4C2:	Data_o <= 8'h03;
				12'h4C3:	Data_o <= 8'hF4;

				// 305 8a1
				12'h4C4:	Data_o <= 8'h00;
				12'h4C5:	Data_o <= 8'hFA;
				12'h4C6:	Data_o <= 8'h04;
				12'h4C7:	Data_o <= 8'h70;

				// 306 1#g1
				12'h4C8:	Data_o <= 8'h07;
				12'h4C9:	Data_o <= 8'hD0;
				12'h4CA:	Data_o <= 8'h04;
				12'h4CB:	Data_o <= 8'hB3;

				// 307 4f1
				12'h4CC:	Data_o <= 8'h01;
				12'h4CD:	Data_o <= 8'hF4;
				12'h4CE:	Data_o <= 8'h05;
				12'h4CF:	Data_o <= 8'h97;

				// 308 4f1
				12'h4D0:	Data_o <= 8'h01;
				12'h4D1:	Data_o <= 8'hF4;
				12'h4D2:	Data_o <= 8'h05;
				12'h4D3:	Data_o <= 8'h97;

				// 309 8e1
				12'h4D4:	Data_o <= 8'h00;
				12'h4D5:	Data_o <= 8'hFA;
				12'h4D6:	Data_o <= 8'h05;
				12'h4D7:	Data_o <= 8'hEC;

				// 310 1e1
				12'h4D8:	Data_o <= 8'h07;
				12'h4D9:	Data_o <= 8'hD0;
				12'h4DA:	Data_o <= 8'h05;
				12'h4DB:	Data_o <= 8'hEC;

				// 311 2-
				12'h4DC:	Data_o <= 8'h03;
				12'h4DD:	Data_o <= 8'hE8;
				12'h4DE:	Data_o <= 8'h00;
				12'h4DF:	Data_o <= 8'h00;

				default:	Data_o <= 8'h00;
			endcase
		end
	end

endmodule
`default_nettype wire

