// 230702

`default_nettype none
module Player #(
	parameter  CLOCK_HZ = 10_000_000
)(
	input wire Clock,
	input wire Reset,
	input wire Play_i,
	input wire Stop_i,
	output wire SoundWave_o
);
	
	
	
endmodule
`default_nettype wire
